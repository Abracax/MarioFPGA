//-------------------------------------------------------------------------
//      lab8.sv                                                          --
//      Christine Chen                                                   --
//      Fall 2014                                                        --
//                                                                       --
//      Modified by Po-Han Huang                                         --
//      10/06/2017                                                       --
//                                                                       --
//      Fall 2017 Distribution                                           --
//                                                                       --
//      For use with ECE 385 Lab 8                                       --
//      UIUC ECE Department                                              --
//-------------------------------------------------------------------------
import Numbers::*;

module final_top( input               CLOCK_50,
             input        [3:0]  KEY,          //bit 0 is set up as Reset
             output logic [6:0]  HEX0, HEX1, //HEX2, HEX3, HEX4, HEX5, HEX6, HEX7,
             // VGA Interface 
             output logic [7:0]  VGA_R,        //VGA Red
                                 VGA_G,        //VGA Green
                                 VGA_B,        //VGA Blue
             output logic        VGA_CLK,      //VGA Clock
                                 VGA_SYNC_N,   //VGA Sync signal
                                 VGA_BLANK_N,  //VGA Blank signal
                                 VGA_VS,       //VGA virtical sync signal
                                 VGA_HS,       //VGA horizontal sync signal
             // CY7C67200 Interface
             inout  wire  [15:0] OTG_DATA,     //CY7C67200 Data bus 16 Bits
             output logic [1:0]  OTG_ADDR,     //CY7C67200 Address 2 Bits
             output logic        OTG_CS_N,     //CY7C67200 Chip Select
                                 OTG_RD_N,     //CY7C67200 Write
                                 OTG_WR_N,     //CY7C67200 Read
                                 OTG_RST_N,    //CY7C67200 Reset
             input               OTG_INT,      //CY7C67200 Interrupt
             // SDRAM Interface for Nios II Software
             output logic [12:0] DRAM_ADDR,    //SDRAM Address 13 Bits
             inout  wire  [31:0] DRAM_DQ,      //SDRAM Data 32 Bits
             output logic [1:0]  DRAM_BA,      //SDRAM Bank Address 2 Bits
             output logic [3:0]  DRAM_DQM,     //SDRAM Data Mast 4 Bits
             output logic        DRAM_RAS_N,   //SDRAM Row Address Strobe
                                 DRAM_CAS_N,   //SDRAM Column Address Strobe
                                 DRAM_CKE,     //SDRAM Clock Enable
                                 DRAM_WE_N,    //SDRAM Write Enable
                                 DRAM_CS_N,    //SDRAM Chip Select
                                 DRAM_CLK,      //SDRAM Clock
			output logic   [19:0]		SRAM_ADDR,
            output logic          		SRAM_CE_N,
            inout logic    [15:0]		SRAM_DQ,
            output logic          		SRAM_LB_N,
            output logic          		SRAM_OE_N,
            output logic          		SRAM_UB_N,
            output logic          		SRAM_WE_N
    );
    
    logic Reset_h, Clk, is_ball;
    logic [15:0] keycode;
    logic [9:0] DrawX, DrawY;
    logic [15:0] MarioX = MARIO_X_LEFT;
    logic [15:0] MarioY = MARIO_Y_LEFT;
    logic [15:0] mushX = 16'd480;
    logic [15:0] mushY = GND_HEIGHT - MUSHROOM_Y_SIZE;
    logic [7:0] MarioAlive = 8'd1;
    logic [7:0] mushAlive = 8'd1;
    logic [15:0] X,Y;
    logic [23:0] RGB;
    logic [3:0] Sprite;
    logic [15:0] screen_offset;
	 logic [7:0] marioState;
    
//    logic [3:0] Mario_Animation;


    assign SRAM_CE_N = 1'b0;
    assign SRAM_UB_N = 1'b0;
    assign SRAM_LB_N = 1'b0;
    assign SRAM_OE_N = 1'b0;
    assign SRAM_WE_N = 1'b1;

    assign RGB = {SRAM_DQ[15:11],3'd0,SRAM_DQ[10:6],2'd0,SRAM_DQ[5:0],3'd0}; 
	
    
    assign Clk = CLOCK_50;
    always_ff @ (posedge Clk) begin
        Reset_h <= ~(KEY[0]);        // The push buttons are active low
    end
    
    logic [1:0] hpi_addr;
    logic [15:0] hpi_data_in, hpi_data_out;
    logic hpi_r, hpi_w, hpi_cs, hpi_reset;
	 logic [7:0] scores;
	 
	 assign scores = mushAlive - 8'b1;
    
    // Interface between NIOS II and EZ-OTG chip
    hpi_io_intf hpi_io_inst(
                            .Clk(Clk),
                            .Reset(Reset_h),
                            // signals connected to NIOS II
                            .from_sw_address(hpi_addr),
                            .from_sw_data_in(hpi_data_in),
                            .from_sw_data_out(hpi_data_out),
                            .from_sw_r(hpi_r),
                            .from_sw_w(hpi_w),
                            .from_sw_cs(hpi_cs),
                            .from_sw_reset(hpi_reset),
                            // signals connected to EZ-OTG chip
                            .OTG_DATA(OTG_DATA),    
                            .OTG_ADDR(OTG_ADDR),    
                            .OTG_RD_N(OTG_RD_N),    
                            .OTG_WR_N(OTG_WR_N),    
                            .OTG_CS_N(OTG_CS_N),
                            .OTG_RST_N(OTG_RST_N)
    );
     
     // You need to make sure that the port names here match the ports in Qsys-generated codes.
     lab8_soc nios_system(
                             .clk_clk(Clk),         
                             .reset_reset_n(1'b1),    // Never reset NIOS
                             .sdram_wire_addr(DRAM_ADDR), 
                             .sdram_wire_ba(DRAM_BA),   
                             .sdram_wire_cas_n(DRAM_CAS_N),
                             .sdram_wire_cke(DRAM_CKE),  
                             .sdram_wire_cs_n(DRAM_CS_N), 
                             .sdram_wire_dq(DRAM_DQ),   
                             .sdram_wire_dqm(DRAM_DQM),  
                             .sdram_wire_ras_n(DRAM_RAS_N),
                             .sdram_wire_we_n(DRAM_WE_N), 
                             .sdram_clk_clk(DRAM_CLK),
                             .keycode_export(keycode),  
                             .otg_hpi_address_export(hpi_addr),
                             .otg_hpi_data_in_port(hpi_data_in),
                             .otg_hpi_data_out_port(hpi_data_out),
                             .otg_hpi_cs_export(hpi_cs),
                             .otg_hpi_r_export(hpi_r),
                             .otg_hpi_w_export(hpi_w),
                             .otg_hpi_reset_export(hpi_reset),
                            .mario_x_export(MarioX),
                            .mario_y_export(MarioY),
                            .mush_x_export(mushX),
                            .mush_y_export(mushY),
                            .mario_alive_export(MarioAlive),
                            .mush_alive_export(mushAlive),
                            .screen_offset_export(screen_offset),
										.mario_state_export(marioState)
    );
    
    // Use PLL to generate the 25MHZ VGA_CLK.
    // You will have to generate it on your own in simulation.
    vga_clk vga_clk_instance(.inclk0(Clk), .c0(VGA_CLK));
    
    // TODO: Fill in the connections for the rest of the modules 
    VGA_controller vga_controller_instance(.Reset(Reset_h), .*);  
								
								
    // Which signal should be frame_clk?
    // ball ball_instance(
	// 			 .Clk,                // 50 MHz clock
	// 			 .Reset(Reset_h),              // Active-high reset signal
	// 			 .frame_clk(VGA_VS),          // The clock indicating a new frame (~60Hz)
	// 			 .*
	//  );

    mario mario_instance(
				 .Clk,                // 50 MHz clock
				 .Reset(Reset_h),              // Active-high reset signal
				 .frame_clk(VGA_VS),          // The clock indicating a new frame (~60Hz)
	 );
	 
    // readRAM marioRAM(.Addr(SRAM_ADDR),.*);
    color_mapper color_instance(.Data_In(RGB),.Addr(SRAM_ADDR),.Reset(Reset_h), .Mario_Animation(marioState[3:0]), .*);
    
    // Display keycode on hex display
	 // mogai
    HexDriver hex_inst_0 (scores[3:0], HEX0);
    HexDriver hex_inst_1 (scores[7:4], HEX1);
//	 HexDriver hex_inst_2 (keycode[11:8], HEX2);
//    HexDriver hex_inst_3 (keycode[15:12], HEX3);
//    HexDriver hex_inst_4 (marioState[3:0], HEX4);
//    HexDriver hex_inst_5 (marioState[7:4], HEX5);
//    HexDriver hex_inst_6 (MarioX[9:8], HEX6);
//	 HexDriver hex_inst_7 (MarioX[15:12], HEX7);
//	 HexDriver hex_inst_4 (MarioX[19:16], HEX4);
//    HexDriver hex_inst_5 (MarioX[23:20], HEX5);
//    HexDriver hex_inst_6 (MarioX[27:24], HEX6);
//	 HexDriver hex_inst_7 (MarioX[31:28], HEX7);
//    HexDriver hex_inst_5 (MarioY[7:4], HEX5);
//	 HexDriver hex_inst_6 (Sprite, HEX6);
//    HexDriver hex_inst_1 (RGB[7:4], HEX1  );
//    HexDriver hex_inst_2 (RGB[11:8], HEX2);
//    HexDriver hex_inst_3 (RGB[15:12], HEX3);
//    HexDriver hex_inst_4 (RGB[19:16], HEX4);
//    HexDriver hex_inst_5 (RGB[23:20], HEX5);


endmodule
